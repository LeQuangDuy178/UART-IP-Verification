package vip_pkg;

  import uart_pkg::*;
  import ahb_pkg::*;

endpackage
