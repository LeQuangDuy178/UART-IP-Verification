interface interrupt_if();

  logic interrupt;

endinterface
