package uart_register_pkg;

  import uvm_pkg::*;

  `include "uart_MDR_reg.sv"
  `include "uart_DLL_reg.sv"
  `include "uart_DLH_reg.sv"
  `include "uart_LCR_reg.sv"
  `include "uart_IER_reg.sv"
  `include "uart_FSR_reg.sv"
  `include "uart_TBR_reg.sv"
  `include "uart_RBR_reg.sv"

endpackage
